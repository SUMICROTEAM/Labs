--------------------------------------------------------------------------------
--
-- LAB #3
--
--------------------------------------------------------------------------------

Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity bitstorage is
	port(bitin: in std_logic;
		 enout: in std_logic;
		 writein: in std_logic;
		 bitout: out std_logic);
end entity bitstorage;

architecture memlike of bitstorage is
	signal q: std_logic := '0';
begin
	process(writein) is
	begin
		if (rising_edge(writein)) then
			q <= bitin;
		end if;
	end process;
	
	-- Note that data is output only when enout = 0	
	bitout <= q when enout = '0' else 'Z';
end architecture memlike;

--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity fulladder is
    port (a : in std_logic;
          b : in std_logic;
          cin : in std_logic;
          sum : out std_logic;
          carry : out std_logic
         );
end fulladder;

architecture addlike of fulladder is
begin
  sum   <= a xor b xor cin; 
  carry <= (a and b) or (a and cin) or (b and cin); 
end architecture addlike;


--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity register8 is
	port(datain: in std_logic_vector(7 downto 0);
	     enout:  in std_logic;
	     writein: in std_logic;
	     dataout: out std_logic_vector(7 downto 0));
end entity register8;

architecture memmy of register8 is

	component bitstorage
		port(bitin: in std_logic;
		 	 enout: in std_logic;
		 	 writein: in std_logic;
		 	 bitout: out std_logic);
	end component;
	
	signal i: integer RANGE 0 to 7 := 0;
	
begin

GenCommand:	for i in 0 to 7 generate
		Li: bitstorage port map (datain(i),enout,writein,dataout(i));
	end generate;
	
end architecture memmy;

--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity register32 is
	port(datain: in std_logic_vector(31 downto 0);
		 enout32,enout16,enout8: in std_logic;
		 writein32, writein16, writein8: in std_logic;
		 dataout: out std_logic_vector(31 downto 0));
end entity register32;

architecture biggermem of register32 is
	component register8 
		port(datain: in std_logic_vector(7 downto 0);
			enout:  in std_logic;
			writein: in std_logic;
			dataout: out std_logic_vector(7 downto 0));
	end component register8; 
	signal en8,en16,en32: std_logic := '1';
	signal write8,write16,write32: std_logic := '0';
begin

	en32 <= enout32;
	en16 <= enout32 AND enout16;
	en8 <= enout32 AND enout16 AND enout8;

	write32 <= writein32;
	write16 <= writein32 OR writein16;
	write8 <= writein32 OR writein16 OR writein8;


	B1: register8 port map (datain(7 downto 0),en8,write8,dataout(7 downto 0));
	B2: register8 port map (datain(15 downto 8),en16,write16,dataout(15 downto 8));
	B3: register8 port map (datain(23 downto 16),en32,write32,dataout(23 downto 16));
	B4: register8 port map (datain(31 downto 24),en32,write32,dataout(31 downto 24));
end architecture biggermem;

--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity adder_subtracter is
	port(	datain_a: in std_logic_vector(31 downto 0);
		datain_b: in std_logic_vector(31 downto 0);
		add_sub: in std_logic;
		dataout: out std_logic_vector(31 downto 0);
		co: out std_logic);
end entity adder_subtracter;

architecture calc of adder_subtracter is
	component fulladder
		port (a : in std_logic;
			  b : in std_logic;
			  cin : in std_logic;
			  sum : out std_logic;
			  carry : out std_logic
			 );
	end component fulladder;
	
	signal cout: std_logic_vector(31 downto 0);
	signal i: integer range 0 to 31 := 0;
	signal Bdata: std_logic_vector(31 downto 0);
	
begin

	with add_sub select
	Bdata <= NOT datain_b when '1',
			datain_b when '0',
			"XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX" when others;

		B0: fulladder port map (datain_a(0),Bdata(0),add_sub,dataout(0),cout(0));
L1:	for i in 1 to 31 generate
		Bi: fulladder port map (datain_a(i),Bdata(i),cout(i-1),dataout(i),cout(i));
	end generate;

	co <= cout(31);
	
end architecture calc;

--------------------------------------------------------------------------------
Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity shift_register is
	port(	datain: in std_logic_vector(31 downto 0);
	   	dir: in std_logic;
		shamt:	in std_logic_vector(4 downto 0);
		dataout: out std_logic_vector(31 downto 0));
end entity shift_register;

architecture shifter of shift_register is

SIGNAL inputs: std_logic_vector(5 downto 0);

begin

inputs <= dir & shamt;
with inputs select 
	dataout(31 downto 0) <= datain(30 downto 0) & '0' when "000001",
		  	        datain(29 downto 0) & '0' & '0' when "000010",
				datain(28 downto 0) & '0' & '0' & '0' when "000011",
		  	       '0' & datain(31 downto 1) when "100001",
		  	       '0' & '0' & datain(31 downto 2) when "100010",
			       '0' & '0' & '0' & datain(31 downto 3) when "100011",
		   	       datain(31 downto 0) when others;
		
end architecture shifter;  



